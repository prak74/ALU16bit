entity Testbench is
end Testbench;
architecture tb of Testbench is
	signal A, B  : bit_vector(15 downto 0); -- ALU-inputs
	signal s0,s1 : bit; --additional inputs
	signal R 	 : bit_vector(15 downto 0); -- final bit_vector output
	signal c_out, z_out : bit;-- final bit outputs
	signal actual_output : bit_vector(15 downto 0); --for checking
	
	component ALU_16 is
		port(
		A,B    : in bit_vector(15 downto 0);
		S0, S1 : in bit;
		R      : out bit_vector(15 downto 0);
		c,z    : out bit
			  );
	end component;
	
begin
-- Connecting test bench signals with ALU.vhd
dut_instance: ALU_16
port map (S0 => s0, S1 => s1, A => A, B => B, R => R, z => z_out, c => c_out);
process-- inputs
	begin
		A <= "0000000000000000"; -- 0
		B <= "0000000000000000"; -- 0
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "0000000000000000"; -- 0
		B <= "0000000000000000"; -- 0
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "0000000000000000"; -- 0
		B <= "0000000000000000"; -- 0
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111111111111"; -- -1
		wait for 5ns;

		A <= "0000000000000000"; -- 0
		B <= "0000000000000000"; -- 0
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "1111001010011011"; -- -3429
		B <= "0000010100001101"; -- 1293
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1111011110101000"; -- -2136
		wait for 5ns;

		A <= "1111001010011011"; -- -3429
		B <= "0000010100001101"; -- 1293
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1110110110001110"; -- -4722
		wait for 5ns;

		A <= "1111001010011011"; -- -3429
		B <= "0000010100001101"; -- 1293
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111111110110"; -- -10
		wait for 5ns;

		A <= "1111001010011011"; -- -3429
		B <= "0000010100001101"; -- 1293
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1111011110010110"; -- -2154
		wait for 5ns;

		A <= "1001001010101011"; -- -27989
		B <= "0010011110011001"; -- 10137
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1011101001000100"; -- -17852
		wait for 5ns;

		A <= "1001001010101011"; -- -27989
		B <= "0010011110011001"; -- 10137
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0110101100010010"; -- -38126
		wait for 5ns;

		A <= "1001001010101011"; -- -27989
		B <= "0010011110011001"; -- 10137
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111110101110110"; -- -650
		wait for 5ns;

		A <= "1001001010101011"; -- -27989
		B <= "0010011110011001"; -- 10137
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1011010100110010"; -- -19150
		wait for 5ns;

		A <= "0111001010100000"; -- 29344
		B <= "0111011110100111"; -- 30631
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1110101001000111"; -- 59975
		wait for 5ns;

		A <= "0111001010100000"; -- 29344
		B <= "0111011110100111"; -- 30631
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1111101011111001"; -- -1287
		wait for 5ns;

		A <= "0111001010100000"; -- 29344
		B <= "0111011110100111"; -- 30631
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1000110101011111"; -- -29345
		wait for 5ns;

		A <= "0111001010100000"; -- 29344
		B <= "0111011110100111"; -- 30631
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0000010100000111"; -- 1287
		wait for 5ns;

		A <= "0111100110000101"; -- 31109
		B <= "0100000001111100"; -- 16508
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1011101000000001"; -- 47617
		wait for 5ns;

		A <= "0111100110000101"; -- 31109
		B <= "0100000001111100"; -- 16508
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0011100100001001"; -- 14601
		wait for 5ns;

		A <= "0111100110000101"; -- 31109
		B <= "0100000001111100"; -- 16508
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1011111111111011"; -- -16389
		wait for 5ns;

		A <= "0111100110000101"; -- 31109
		B <= "0100000001111100"; -- 16508
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0011100111111001"; -- 14841
		wait for 5ns;

		A <= "1110101001001001"; -- -5559
		B <= "1101101000001011"; -- -9717
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1100010001010100"; -- -15276
		wait for 5ns;

		A <= "1110101001001001"; -- -5559
		B <= "1101101000001011"; -- -9717
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0001000000111110"; -- 4158
		wait for 5ns;

		A <= "1110101001001001"; -- -5559
		B <= "1101101000001011"; -- -9717
		s0 <= '0';
		s1 <= '1';
		actual_output <= "0011010111110110"; -- 13814
		wait for 5ns;

		A <= "1110101001001001"; -- -5559
		B <= "1101101000001011"; -- -9717
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0011000001000010"; -- 12354
		wait for 5ns;

		A <= "0001011000111011"; -- 5691
		B <= "0110100011101110"; -- 26862
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0111111100101001"; -- 32553
		wait for 5ns;

		A <= "0001011000111011"; -- 5691
		B <= "0110100011101110"; -- 26862
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1010110101001101"; -- -21171
		wait for 5ns;

		A <= "0001011000111011"; -- 5691
		B <= "0110100011101110"; -- 26862
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111111010101"; -- -43
		wait for 5ns;

		A <= "0001011000111011"; -- 5691
		B <= "0110100011101110"; -- 26862
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0111111011010101"; -- 32469
		wait for 5ns;

		A <= "0000001010010010"; -- 658
		B <= "0100010111001000"; -- 17864
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0100100001011010"; -- 18522
		wait for 5ns;

		A <= "0000001010010010"; -- 658
		B <= "0100010111001000"; -- 17864
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1011110011001010"; -- -17206
		wait for 5ns;

		A <= "0000001010010010"; -- 658
		B <= "0100010111001000"; -- 17864
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111101111111"; -- -129
		wait for 5ns;

		A <= "0000001010010010"; -- 658
		B <= "0100010111001000"; -- 17864
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0100011101011010"; -- 18266
		wait for 5ns;

		A <= "0110111001101010"; -- 28266
		B <= "1100001101000100"; -- -15548
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0011000110101110"; -- 12718
		wait for 5ns;

		A <= "0110111001101010"; -- 28266
		B <= "1100001101000100"; -- -15548
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1010101100100110"; -- 43814
		wait for 5ns;

		A <= "0110111001101010"; -- 28266
		B <= "1100001101000100"; -- -15548
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1011110110111111"; -- -16961
		wait for 5ns;

		A <= "0110111001101010"; -- 28266
		B <= "1100001101000100"; -- -15548
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1010110100101110"; -- -21202
		wait for 5ns;

		A <= "1110101001010100"; -- -5548
		B <= "0001010110101100"; -- 5548
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "1110101001010100"; -- -5548
		B <= "0001010110101100"; -- 5548
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1101010010101000"; -- -11096
		wait for 5ns;

		A <= "1110101001010100"; -- -5548
		B <= "0001010110101100"; -- 5548
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111111111011"; -- -5
		wait for 5ns;

		A <= "1110101001010100"; -- -5548
		B <= "0001010110101100"; -- 5548
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1111111111111000"; -- -8
		wait for 5ns;

		A <= "1101000000101110"; -- -12242
		B <= "1010000100100001"; -- -24287
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0111000101001111"; -- -36529
		wait for 5ns;

		A <= "1101000000101110"; -- -12242
		B <= "1010000100100001"; -- -24287
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0010111100001101"; -- 12045
		wait for 5ns;

		A <= "1101000000101110"; -- -12242
		B <= "1010000100100001"; -- -24287
		s0 <= '0';
		s1 <= '1';
		actual_output <= "0111111111011111"; -- 32735
		wait for 5ns;

		A <= "1101000000101110"; -- -12242
		B <= "1010000100100001"; -- -24287
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0111000100001111"; -- 28943
		wait for 5ns;

		A <= "1101010100010110"; -- -10986
		B <= "0011010001110101"; -- 13429
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0000100110001011"; -- 2443
		wait for 5ns;

		A <= "1101010100010110"; -- -10986
		B <= "0011010001110101"; -- 13429
		s0 <= '1';
		s1 <= '0';
		actual_output <= "1010000010100001"; -- -24415
		wait for 5ns;

		A <= "1101010100010110"; -- -10986
		B <= "0011010001110101"; -- 13429
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1110101111101011"; -- -5141
		wait for 5ns;

		A <= "1101010100010110"; -- -10986
		B <= "0011010001110101"; -- 13429
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1110000101100011"; -- -7837
		wait for 5ns;

		A <= "1001111101011010"; -- -24742
		B <= "0110111001000001"; -- 28225
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0000110110011011"; -- 3483
		wait for 5ns;

		A <= "1001111101011010"; -- -24742
		B <= "0110111001000001"; -- 28225
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0011000100011001"; -- -52967
		wait for 5ns;

		A <= "1001111101011010"; -- -24742
		B <= "0110111001000001"; -- 28225
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111000110111111"; -- -3649
		wait for 5ns;

		A <= "1001111101011010"; -- -24742
		B <= "0110111001000001"; -- 28225
		s0 <= '1';
		s1 <= '1';
		actual_output <= "1111000100011011"; -- -3813
		wait for 5ns;

		A <= "1111111111111111"; -- 65535
		B <= "1111111111111111"; -- 65535
		s0 <= '0';
		s1 <= '0';
		actual_output <= "1111111111111110"; -- -2
		wait for 5ns;

		A <= "1111111111111111"; -- 65535
		B <= "1111111111111111"; -- 65535
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "1111111111111111"; -- 65535
		B <= "1111111111111111"; -- 65535
		s0 <= '0';
		s1 <= '1';
		actual_output <= "0000000000000000"; -- -65536
		wait for 5ns;

		A <= "1111111111111111"; -- 65535
		B <= "1111111111111111"; -- 65535
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "0000000000000001"; -- 1
		B <= "0000000000000001"; -- 1
		s0 <= '0';
		s1 <= '0';
		actual_output <= "0000000000000010"; -- 2
		wait for 5ns;

		A <= "0000000000000001"; -- 1
		B <= "0000000000000001"; -- 1
		s0 <= '1';
		s1 <= '0';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

		A <= "0000000000000001"; -- 1
		B <= "0000000000000001"; -- 1
		s0 <= '0';
		s1 <= '1';
		actual_output <= "1111111111111110"; -- -2
		wait for 5ns;

		A <= "0000000000000001"; -- 1
		B <= "0000000000000001"; -- 1
		s0 <= '1';
		s1 <= '1';
		actual_output <= "0000000000000000"; -- 0
		wait for 5ns;

end process;
end tb ;